module segmen7(m,HEX0);

	input [3:0]m;
	output [6:0]HEX0;
	
	assign HEX0 = 	(m[3:0] == 4'b0000)? 7'b1000000 :	//0
						(m[3:0] == 4'b0001)? 7'b1111001 :	//1
						(m[3:0] == 4'b0010)? 7'b0100100 :	//2
						(m[3:0] == 4'b0011)? 7'b0011000 :	//3
						(m[3:0] == 4'b0100)? 7'b0011001 :	//4
						(m[3:0] == 4'b0101)? 7'b0010010 :	//5
						(m[3:0] == 4'b0110)? 7'b0000010 :	//6
						(m[3:0] == 4'b0111)? 7'b1110000 :	//7
						(m[3:0] == 4'b1000)? 7'b0000000 : 	//8
						(m[3:0] == 4'b1001)? 7'b0010000 : 7'b0111111 ; //9
			 
endmodule