module lab2part1(SW,HEX0,HEX1,HEX2,HEX3);

	input [15:0]SW;
	output [6:0]HEX0,HEX1,HEX2,HEX3;
	
	assign HEX0 = 	(SW[3:0]==4'b0000)? 7'b1000000 :
						(SW[3:0]==4'b0001)? 7'b1111001 :
						(SW[3:0]==4'b0010)? 7'b0100100 :
						(SW[3:0]==4'b0011)? 7'b0110000 :
						(SW[3:0]==4'b0100)? 7'b0011001 :
						(SW[3:0]==4'b0101)? 7'b0010010 :
						(SW[3:0]==4'b0110)? 7'b0000010 :
						(SW[3:0]==4'b0111)? 7'b1111000 :
						(SW[3:0]==4'b1000)? 7'b0000000 :
						(SW[3:0]==4'b1001)? 7'b0011000 : 7'b0111111;
		
	assign HEX1 = 	(SW[7:4]==4'b0000)? 7'b1000000 :
						(SW[7:4]==4'b0001)? 7'b1111001 :
						(SW[7:4]==4'b0010)? 7'b0100100 :
						(SW[7:4]==4'b0011)? 7'b0110000 :
						(SW[7:4]==4'b0100)? 7'b0011001 :
						(SW[7:4]==4'b0101)? 7'b0010010 :
						(SW[7:4]==4'b0110)? 7'b0000010 :
						(SW[7:4]==4'b0111)? 7'b1111000 :
						(SW[7:4]==4'b1000)? 7'b0000000 :
						(SW[7:4]==4'b1001)? 7'b0011000 : 7'b0111111;
						
	assign HEX2 = 	(SW[11:8]==4'b0000)? 7'b1000000 :
						(SW[11:8]==4'b0001)? 7'b1111001 :
						(SW[11:8]==4'b0010)? 7'b0100100 :
						(SW[11:8]==4'b0011)? 7'b0110000 :
						(SW[11:8]==4'b0100)? 7'b0011001 :
						(SW[11:8]==4'b0101)? 7'b0010010 :
						(SW[11:8]==4'b0110)? 7'b0000010 :
						(SW[11:8]==4'b0111)? 7'b1111000 :
						(SW[11:8]==4'b1000)? 7'b0000000 :
						(SW[11:8]==4'b1001)? 7'b0011000 : 7'b0111111;
						
	assign HEX3 = 	(SW[15:12]==4'b0000)? 7'b1000000 :
						(SW[15:12]==4'b0001)? 7'b1111001 :
						(SW[15:12]==4'b0010)? 7'b0100100 :
						(SW[15:12]==4'b0011)? 7'b0110000 :
						(SW[15:12]==4'b0100)? 7'b0011001 :
						(SW[15:12]==4'b0101)? 7'b0010010 :
						(SW[15:12]==4'b0110)? 7'b0000010 :
						(SW[15:12]==4'b0111)? 7'b1111000 :
						(SW[15:12]==4'b1000)? 7'b0000000 :
						(SW[15:12]==4'b1001)? 7'b0011000 : 7'b0111111;
						
endmodule
						