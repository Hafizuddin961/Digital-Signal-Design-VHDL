module comparatorA1(SW,cA1);

	input [15:12]SW;
	output cA1;
	
	assign cA1 = (SW[15:12]>4'd9)? 1:0;

endmodule



module comparatorA0(SW,cA0);

	input [11:8]SW;
	output cA0;
	
	assign cA0 = (SW[11:8]>4'd9)? 1:0;

endmodule



module A1segmen7(SW,HEX7);

	input [15:12]SW;
	output [6:0]HEX7;
	
	assign HEX7 = 	(SW[15:12] == 4'b0000)? 7'b1000000 :	//0
						(SW[15:12] == 4'b0001)? 7'b1111001 :	//1
						(SW[15:12] == 4'b0010)? 7'b0100100 :	//2
						(SW[15:12] == 4'b0011)? 7'b0011000 :	//3
						(SW[15:12] == 4'b0100)? 7'b0011001 :	//4
						(SW[15:12] == 4'b0101)? 7'b0010010 :	//5
						(SW[15:12] == 4'b0110)? 7'b0000010 :	//6
						(SW[15:12] == 4'b0111)? 7'b1110000 :	//7
						(SW[15:12] == 4'b1000)? 7'b0000000 : 	//8
						(SW[15:12] == 4'b1001)? 7'b0010000 : 7'b0111111 ; //9
			 
endmodule



module A0segmen7(SW,HEX6);

	input [11:8]SW;
	output [6:0]HEX6;
	
	assign HEX6 = 	(SW[11:8] == 4'b0000)? 7'b1000000 :	//0
						(SW[11:8] == 4'b0001)? 7'b1111001 :	//1
						(SW[11:8] == 4'b0010)? 7'b0100100 :	//2
						(SW[11:8] == 4'b0011)? 7'b0011000 :	//3
						(SW[11:8] == 4'b0100)? 7'b0011001 :	//4
						(SW[11:8] == 4'b0101)? 7'b0010010 :	//5
						(SW[11:8] == 4'b0110)? 7'b0000010 :	//6
						(SW[11:8] == 4'b0111)? 7'b1110000 :	//7
						(SW[11:8] == 4'b1000)? 7'b0000000 : //8
						(SW[11:8] == 4'b1001)? 7'b0010000 : 7'b0111111 ; //9
			 
endmodule