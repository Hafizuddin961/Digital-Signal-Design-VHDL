module comparatorB1(SW,cB1);

	input [7:4]SW;
	output cB1;
	
	assign cB1 = (SW[7:4]>4'd9)? 1:0;

endmodule



module comparatorB0(SW,cB0);

	input [3:0]SW;
	output cB0;
	
	assign cB0 = (SW[3:0]>4'd9)? 1:0;

endmodule



module B1segmen7(SW,HEX5);

	input [7:4]SW;
	output [6:0]HEX5;
	
	assign HEX5 = 	(SW[7:4] == 4'b0000)? 7'b1000000 :	//0
						(SW[7:4] == 4'b0001)? 7'b1111001 :	//1
						(SW[7:4] == 4'b0010)? 7'b0100100 :	//2
						(SW[7:4] == 4'b0011)? 7'b0011000 :	//3
						(SW[7:4] == 4'b0100)? 7'b0011001 :	//4
						(SW[7:4] == 4'b0101)? 7'b0010010 :	//5
						(SW[7:4] == 4'b0110)? 7'b0000010 :	//6
						(SW[7:4] == 4'b0111)? 7'b1110000 :	//7
						(SW[7:4] == 4'b1000)? 7'b0000000 : 	//8
						(SW[7:4] == 4'b1001)? 7'b0010000 : 7'b0111111 ; //9
			 
endmodule



module B0segmen7(SW,HEX4);

	input [3:0]SW;
	output [6:0]HEX4;
	
	assign HEX4 = 	(SW[3:0] == 4'b0000)? 7'b1000000 :	//0
						(SW[3:0] == 4'b0001)? 7'b1111001 :	//1
						(SW[3:0] == 4'b0010)? 7'b0100100 :	//2
						(SW[3:0] == 4'b0011)? 7'b0011000 :	//3
						(SW[3:0] == 4'b0100)? 7'b0011001 :	//4
						(SW[3:0] == 4'b0101)? 7'b0010010 :	//5
						(SW[3:0] == 4'b0110)? 7'b0000010 :	//6
						(SW[3:0] == 4'b0111)? 7'b1110000 :	//7
						(SW[3:0] == 4'b1000)? 7'b0000000 :  //8
						(SW[3:0] == 4'b1001)? 7'b0010000 : 7'b0111111 ; //9
			 
endmodule